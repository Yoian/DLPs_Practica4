
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Ejercicio4 is
end Ejercicio4;

architecture Behavioral of Ejercicio4 is

begin


end Behavioral;

